defparam AESL_inst_MultipleToSerial.tmp_elements_num_loc_channel_U.DEPTH = 11'd1000;
defparam AESL_inst_MultipleToSerial.tmp_elements_num_loc_channel_U.ADDR_WIDTH = 32'd10;
